BZh91AY&SY�R� �߀Py���w߰����`�< �p0�� @
 ( �� ��z�� d   ��5O�7���@�4 h � hT��EI�       �mS=S�ɣ 4     4MR�h P      D� )�)��4MCz�4y�=&�U?@	T�&L�  @a107�5�+��AS@1>$U�>_��?27�#	n�Q0?H]RP�Eo���J��f�0;v����.�޻;::;I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$���tua���뤒I$�I$�I$�I$�I$�I$�I$�I$�I$�I&8���ɥ��_f��1���,϶yB�h�-y��{� ���{��#���*SF�P�]��"4��e`ҳ�B��l�;�[���i�\�;5]��ц�R��St�]Y�����$2�w��}~bv�m��yk�e��Ûp�ױ�L�8#��S��]dγ��{�]�\P�-eG�M���P��oBIŊ#�����5�<4�˛T�k���r�^R���b��������λ���p<�*�����Aj.�v]&nQ��7b�z��+�Y�
�m�xC<��F��ܳ���|����]z5�"e|:7������&�V�pJ�(K����m�����|�f��[G�nW,�5�}�9��T{B�R�IgY�P�*dV�*_l+��W=��x����]��Y��٫n�@9+ϰ��>�������k�H _ğ�1���g�N_��������(��,�c��I$�I$�I$�I$�I$�I$�I$�I$�L��Ƽi�1�6d�3f͚I$�I$�I$�I$�I$�I$�I$�I$�8a:�Qyp����ȷ��U�ͤ�Q�u`���ڨj�]�\���0*!ei��ʫI&sB�E�QT��u�B�3]d+��C8-B��^	�D�:��v7�~fUwo�<���X��N����.��ȣy��p9���A�	�yU����4w�_�����fku��C�4@�2�(��,Gؾ�w�:�7߳��4��1��iƇ��n��P�Ac0�D������a�D�\�'�8ߴ��
�x���h!��y4�4Z3�V���������1��G"Xӝ}�Um�E���0"�'	�Z.(iq5�����I�x�
�����B�"&�S�t`�n�)���C�V�ݡp~����9�]�Sf���o��cOq�K,��,�ΨgRC�<(#D��_/�_0�����������LE@%�0x��<!���_�"�|�Q?tk�P�����"��A�`������3���7F(@hxo��ǆ=��$���L�$#�G���<#�(�.�q	 �C!�?�aU�o�~0bDH��Ŋb�K�x\J*u����!A�2�a���N�;�K+(� ���q��i��hq/,N�s��i�ꭣ��x�F�_;�ˎ��J�_3��b��<U���,��9%�/�6�Ӵ?谡�X�hHq�Cn�!��T���G=(��	>rG	�cH,��<A:̀�P�}�Ae��'L��D8���xh2�3�;�4}�q�8����q�V}��F��3�(�=�iC}�$�<9��4�qg� D������{��"	�I4�0���=/��ɽ�޳�mW*�>�{o�M^��ʯT���G�4��30�0³Q�I!�����Gؖ�4�9#�<bTqG�(a�=���E�&!�4bg�Nzj
���G�I(�H�OB��dT3x�0Rt"�aݨ$��x��Ǌ2���'��ؠ�N(��x�8W摙��I�9�l�@���j(�T1h��Y��Ë���`�H�����wf��h��=�3��I���e��(ľ�È���<Yƚl�~��';S~�5$ь�Y���ٵ��d|�7�ƈ�U�L��Q�a�va�a�O�#P���4f�t`�A�A�,sG��ʽ�����$b�sKᰂ%-)\��8-H�Q��cw�3Pp��Y���(��!���a|�q�WIh����,�����IQ��_"K��$@W%c�p�(6�4~ o�1�ǆjI
�90!qP`�hP}'y*N��7(�(,�,�=�yP�[�\D�0xC�W{U!âOA�Oi�����㫙A��˻��h��9t�0jd���H��*]4#'�N�Z��mI,XŒaƛ�a�a'�Lt3&��1�C�x�DYf�*��!�~����Ēp�g��G6	+�>J�,��5"��1��(�H04���Ƣ~�� �K�ϑ&A�_1L�1_���8��$��AL��~`����$��L�������a����$8��`<� o�,���0��A�!��Qĕ#�r�	$��<g��d[d5`�6[���=���C�:CO�5Vg�UA=^�w/���MƐi�ie�Ye�Y��G�ID��6�;Ry$�q:J��C`X8�P�1�I��;5|i���,��,aI3S�����9P�G��0��N���#H4ӏ?Ne�Q�S���9~<1�|�S� ��.�K��0���aGL�35��J�#�9�B/�o.�a��|�z�}eN��ؒ�fV}�����K+�*"�Pi��C�h�=j����8��۵��՛��Mx��ڳb5}ZpŒQF�a�a���.u�����=�AÞ�E��?}�I+���e8�r�O���,҆�$�	ɉ��!ڏ�����@�0���
as�aC(,<0�l��Bwj����q��Fy4b<1��5ADr��}�$�G8�����T>��|b�G�¼a��fg��8�|��G��{N�8��<�f��/�gO6��u
^���'^����++���A��<Њ��<G�lE��k�!~$�KÌp�"���P�bа�ȹ*ؓ�1���	\�E&'�Bh���?E� ��^"E�C�(���A.�h�X��i9�|�G��� �2ؑ0b�1?H�M�b����E��#9B�M�������h��.T��1���Ѵ�J
'֚U�}�g1����#K<i�,K�.�h#s�MT�5�&F��]�&8��	�B7��}�tQ��r)�����C�4��9e�Y��ҹ��3.4G�����8�Otc��:(>��qQƖA1��Gǈ(m�c�^d<�i ф9#�0�k�H�IE��zS��3C�01#y{��4�/�8��hQ�<�h�,A%��'�)��f��8�L8��E�gG�p^�&#��z�@�'������+I%x�UU5��q��;o?�=#����������*��6Iq�D��Ak�q�p�%#��䒖�RDL�M������?nJ^3ޝ���n��	�h�MD"h���3��&��4B&��7:t1D��D"h�Mrg,D��,D���������M�ܛ���4X�D"n��	B[:8��#I��H$�FH�. �gn1#I�	����շL�;��ނ��
o��<�a���"_E��Sx�I��1�i����C#.1��Bl,��P���d�Ǉ��<��!D��d�*����J���DW�&��|}�F�Zz��6Pd'0E}iN� ������������~W�(�
C�Z����5��:�=�"��xO�?]�!x{#lP���o��4斂B%���}_�B�>&9�K���[��<	����Q�}�:�D���PAP��"��n�gXڛ)�����rcI�e2FY2i�2d$R	 cq��E�����Y,Z��E�zz���IH~cJ`
F
�-�ǎ�9�¶��`ãF<Z�� ��&p<����'�W�ݽ("��!I{d�w�;p����x73�lqd3��W>��s��HA��M|��ekz��8�<{� "�\�I�a�2}ڊ�ӖXe�]�)[�"����'7��A��;�V���^O67&ay�\����U���hl�.m����(as�w���Y�٦Q?���rK8�bc�pK�T1����%�;�wxf!:�N "�^и_?hl
���y���R���h�t�I���v0�<��)?�v��2�Y�A�HD>�ڝ@"�Ǎ���_Ӡ�����t���VI��q$e����رJ�Zf����,��@����u��C�=Ak^_�.l^6�GE�"�7X_E!����hm��ٻ=x���G2� �/�?���lպ)�؞!`�wnLཥ��� ��6�%X�:��/4�^NB��̈́<
��^�@ѩ2?���)�����