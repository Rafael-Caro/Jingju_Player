BZh91AY&SY���w �߀Py���w߰����`�< �>p0��( P�*�	 (  ( � �   *�S��� h ɣL��  �O����       $���SG�2h�A��145IP        (@�О�x���P~�hi�jO��	T� %R��0�&�F0�24ͺM7��í �(*`� d'�Ej��y¯����6�H��Z�P�(��\X�H��n#�m܏O��O�wzw^rI$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$����v�m�Md�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�Y�VXM,�3h���ͫ�a�E��+���^�O���^|�w�To
��LH��6�E����U�*�)Rk{$RneK������}uꪘ0������n��.��a\�W��qV
�z�6�r����ޮ�{a��s:�e�|'wR��w/��Ι�o����G��İ�����zM�Q8��0a{�贪T��V��[����rڦʩi��K����꾪��w}�{'G���0�}UK린�FR�[˫�)
o�<�L����L�iuuh�;�>�⇼P���yEJ���
�3W
�hX�5��c6�`��Ħa̗�z�s�y����a�>�2>W�7*gC��ܨ��b���J��ا
���Y4 �v��
��ږQܼ3���]c�+�ɪOVL��?�~@�������|}�� 3�����p�?*�ǹ��3��D�alZ��I$�I$�I$�I$�I$�I$�I$�I$�e�C1�5c�LX����2d�I$�I$�I$�I$�I$�I$�I$�I'8Y;��˨QD]��+-�N�^�@Q����=v�Rx靂T���,&B���Vi�n�K�V�l�NU���b��}D*r��oP���&�X_�&X[��#[��<<6�X����YWhek�7�
�M��q��d�O�����ڭ}���z8^�J�ƹ���ۃ�Ǹi��aEQEX��}��u�o����L,Әb�ď�rq�s!BHq1C�K�:���qFtK��2q�3�7�\aQ�<GCD4��<�i�-��E���i�qgaf��H�#�,iξ�*�ݢ��g�����-4���>>�,�4�N4��9�e�'���E\V]畠��b�j��mQ���#荒�9�]�Sf���E0�<q�K,��,�ΨgRC�<(#D��_`�`�q~_|�(_P��mf'N6Rb*/�a�ČY���J�(_}�#媉��_ℾ��|H��/�� �t�@�}i���1BC�||h�<1�M�'�f�g� qZ8Ġ�qG��w눈��H���A� ��
��|H@��"D�@�,S^H���QS�����
1����'�t�߂YYE�x�>� ӌ$�M4�q/,_y�c>k�8�b<+,C��4�UvW��q�Ú�_0��Yc�q���Ye�Y�$���&�C��v���=�>a�	0��cM��d5�ʃ�0_�ǥ�A'�H�1 �i�q�������M ����N8����q�9e��0�0�T�C������⎓Do�9�dAY�kƂ�r�8�$���%��$�`���IŞ�[ϟ'��/���h�$|,�$��<E�i�K�D���޷ޣ�rV'�����#��[~;8�#�qf�a�aY��$��pO���#�KBp���ƞ1*8�Ŕ0��p��ȓ�13��'=5`�a��$�Q$}��P?Ȳ*	�<A):}�����<a���b�x��b�Pz'QB<i�+�H���$�Ӝ�g D��5P�D�(($4b�������`�H�����m+"��ƌG}���,yJ�(ľ�ÈsL�Ŝi�W�2��ՙ��I4^t]@�ѥ¬\���[��4D��eZ"�8�+�c0�:~I�}�h٣7�zAc�?�^U�*
7�(<H��#�aJZR�;�pZ�̣�:08��:f��!���e�ag�I<7�c�K�2��KExw�g�/��x�*H"�(�J��_�"�+ۆ�A�9��}�<3RHP�Ɂг�� kB��;�P�uH�q�@-qAdaga�Kʇ�r���$�����ڨ�'��0�O���絬�u-�5GU{{M3o�K�Ƭ$��db�l�"_�,�Ne
�@�aƛ�a�a'�Lt3&��1�C�x�DYf�*��!�~C�kIÐq�,h}�$�l�*,���Ԋ��8�	 �Ӈ7�	�4�I.�>D�H1�|�M2d�|xF����N��J�2s����C#l��Nq2K���kG����B'ð��#�E9�����0�����"�<Q"�8��c�V�I��<xߓ�ȶ�j��l��<C5�^�0N��b�1:3�5y[�^2��K��4�,��,��0�H��	!�"k��yI<�I�8�%y܊�!�,c(q��$�ם��4�XƖQ�0�$���gzk���(r#�J�q�˧a���iǊ��2ъ(�)�����>��1�]���1�a_-4��fj
3	*�GsB�_�2�]��Ǌ�����0�=��%�̬�����WBT"
(E8�i�q��y�F.�����CMSN4���5�s�FDb�
���4�0�0�д	s���d�Xő� ��-~hi���%�I_0��(q�{�R}�FAf�0��'�8NLMu9�}��.� a�.���SC��Aa��d�"�Pf6h���*3ɠaG�0�&�(�Y"�D�h�1�86*����Q�CW��4b�,��8Ç��ŗ��8Ǝ#�?x�N4���J�r�<6�萗��ݝ�5���N��cX��++O�a�q�p�B(r�(�y=�y��.�Q��r�/1�x�$G�B(q�B"�bN��$ys�<9��I	�﯆4�W�αx��@�c;�9��	bOŤ箅�ޗ����bDx����#�7݋��guD�H�k�i4F�&�W�뱣��<�S��h��hVR xF��((�ZiV�<I�Ŝp��JO0�,�4'�J}4�ȬNIz��%�83_UA%�ǆ�����O볡�~T�\�q�qƙ"��,��;>�W#��eƈ� �� r�҉�t��gE�b�!�8�� ¦;:(���1��/2S��h���j5פh$���=)�����`������O�p�4(�g4x� ��L�Ŕ�g3R�w&bB��[3���8/E��=B f���yǴ�+I%x�UU5��q������j�̼��NV�	�	����%kx��8�)"JGs��%-$���h�-)d---"&~�8�.��]�Ӯtn㣄�4B&��4M�puқ��4B&�D�4B&���D�4B,D��!u�C��dM���M�Gh��gM"h�N�p�""!��t:h��D�GD$i	l��6H�d��	6��3��$���H�d�A-)% �m�z�ʅ�h�vT��\#��X�+�ِ�>��1~����j��R`ڕr�؟�T/�P0��N8�=?-�'�}�i��`�ELlz���e���݉������"+�SI�y|zM^����j�b'0E|�gN� ��҈�}���!�xp����,���F��؆���R��WR��O�i\��(������%`��	Zp0Og�C�� Id��_�u�Wq�^SI��$]���i�K_@��
����v<��6S5��&)��dɦDɓH$X�����Z�h�3�bD�ZW����y��Ƈ�9D?qE0�
Q�	 ��0߱�A0��Q�tf�{H�1ᓚ^6� ��m��ݶڔ�+SxQ.j�m�NW������3q[�aT2���N{���B��8����9j���ٛy�nÈ��v�t�n������G�Y�E�눪�:�E����>PxC����R�^6.�x�&Aq�����*�M�a��!]�k
�`���Y������xU�U�
'�Q��.)V�=�L!k7�����DV�pN�]��N�&�_xX_�Xj
E�ϑ��<x���iQ{�t)&�iu�l9�� {�'���n�@dYVz�{R���H���`��.������q�=���������HBRUh�_#�V�q����tcd9e�+[�����团�[�[F����Pj#A�v�^̴�d8��S�\o?���FȤW�bw�C�4�be�\�ۘ�]��J�'QA���<0��o���C�����bm	���ܑN$'�-��