BZh91AY&SY���W �߀Py����߰����`��(�����
(�((�ErqE *�I��2��jz�� h bz��~A���	�	�d�� �0L@0	�h�h`bc�0L@0	�h�h`baD3D�56�&�T�'�� �4zm@�b�� #Fɀ�i�� �	�46`�	R�� 
��
f/����A.#
�OH28E"B1V���*&'��(d�� �D؃Q�Lb������cFv��r.)JR��(�)JR����)JR��)*R��)J)JR��(�)JR����)JR��)*R��)J)JR��)HR��)JR��)JR��(�)JR��)*B��)JR��)JR�,X�p*��.B�|����˳�T`7��]���8�U�f{��Ԩs6I����H���^ޢ��j�[�;&�ֳ����v�n�7t^(��)-�nL;���k$�i��(���aeKF�팷$�P���7;-��DЋM����X�x���[7�Onm<E]5179em"���L��I�C��=Ơ^\#*N���]�� �zfb�g��Ӆ�嬶#��Ƅ�Q�wZa-�@m[���6��׵/j7r�܃
�ә�;v�UԲ��n(2o[�&A��l�v�NВm��Q�Zw��E�6NT��T���\4�v�(�9�2�$JD�ڇ9~��6k��-Y*SO����Z�ZֶV��l�kZ�Zֵ����iw��k����B�m��ֵ�n�Zֵ�n-iZֵ�m��٨��O'Y�q�Z-kZֵ�k-kZֵ�k-kZֶ�m�x�N#q����kZֵֶ�kZֵ���+Z���*�Ys6�f���z�Zػ��[BT�,���B��E��� OP+(�5i+:�N_y�n��a<:ϫ�~P6�$ׂ�̂���P�ڥ�8M�S�)�=0�+Q[�&3��'�8�X֚i�L��,�Yw[DCg1���������-��(�J�s|�b%N)��i��ܶw��-�4�����s���2�[Z��j��v�6ꖇt��V�S�u�/1��B�-�S�b�B^CM/���~	`� '��X��M�-X�f�p�ܗ=�����a��[Zi��~7��mJR���LCC���e�?�R:�NT8�ڈB��]"���u-��6ҷ\�׹ܭ�9�e�[�Ud�m��j#�g��#��+Ĵz>�v��	�%�yM�9���P�5��O�-��!���-?	Z2�)��e��!
��	dA�h��}�{u-�]���b�f�W�c��U��-<�,�ʒ�)JR��"".�6�Z�>[�L��]��F�҉=��e����/��R�OuXc�ی�w��VS��9a�q4�8�LK���Sư�a��e�T�\��S�qo�[��C-��G�yԌ��J5-��YL!�m
|}�y'k��z�}��W�=��Z�����K�Ӿ�����ē['Av)��M)JS:�i�Ziݦq�ȇ���K�RזXT��J}	Nc����Tޣ[�)��|�e�ͥ�<i)�����䶆Py�J(y)u�ؤS(S�n&�j�٘z4����iNe/q�KI1�e!�"��)B� t;�k��(�.]$8��8r�!�g���]T_m�V�Ye�)JR��Z�1�'#��!�]k�q�^wS���e2�_4���f���O�=��
o��b���؋�\3UZ01!d�S�=l�#S�3�\]���wkU�|ӈCi}��8��,�-�Y�Y!�q�e��Լ��mt�O��9��I_VM�4��7�[���]ޭT+2�&�Cۡ���X[��`��?V��)JS����jR�֡����e��y}�#,�#�������:F)m�a��)|���ȧ>��iZDyN=��4��~��Mg/�Qž��}����j�qF�i+|۵9b�������Sv��\�}�E�g\滞�Us�.4�-�9��� ����[�=�4�L�M4�Ye�[�m��P��ji�mM���y��gZ~S�Cf�w�)=\�Xw�v_<�\��o���1�b޴�_>���x�<ϣ�O1�6�km�b+8m�:Ӻ�&�L�msx4�<R��T�iJ��qb�("D��,��4�M5�n&9��R�I}�Z�8���>6�����5�^[�e�9�������H���^�G��Z���u�}�t�~q�K�^m�#=�4ź�|C�Tu,����2�̹��n!�o|���<=g=m�� \���!.(�WE�E(ɔ�4<�[���i��R��Ye�V����~V��hQ%��T���s��1Ō���� D��Ӯ�g����'�Nk���_!�_ᶐ�-I_��<iN%zoDo�|�g��4��ܶ�+C|���Z]���`󜐦r�����K,\Q��Zkuϝeo5��i���*R��p�x�#��
�Jߢgzmxg��F�}�(�X���}U3f[{,���>q�Ԇ��v+�z���b)1�:�9ǖ�=��3o��b>��o�GT٨����Ӵ��!	7�$�A���S�:�^+�Y|�^���_�&�ۘ�&�,�m���4��	b1�	 A�1�v�X�	b0�hS0�X�����`�2%�H�"a��H� @�@� C$� ��Z(
(�
��-�d h��"e<b�Yع�0Ƅ��(�!'|P�P�"뢹����*���妿��*Qw������~5�vVcAhL�ˆ�K�����š��By''h~y�*��5P~��O�@#��뛄�܍܀�����@@OE�h|�c�C���q��޶0B��kG���Csӱ��:{�3�C�>㞟ˬ��R�0X�g�6j@�H��FK�𐢏���Iu�0�'q���<��[X�*5"��ㆹ�K�CB�(��o;X �a��B+� �"�, �0G����idР�x>ڹ ���Y]�A��@� �1��Ko2�t��Xe�mw���|�=-Gpf�ju�F�~z��ׇ���9��D��).�/�GkZ](�Z�mc�GAh�$�=}`������ΰ�|^`�zS�������c��:�4r�g ��##��+�S�n.�<LV!��(�px�|��/�bz�z�M��7Y���0	�,/�m�0���B��[u�F�4D�������� Y�j�fQ?�N.kg<X@��R��A�2��'8�j�WN ���`\��n���=هǭ��F�'����Y�Gk��=L>��EaI��?c���耒��>+��ʍ��F�f���	l�R���������D�r\��.��M\ J�B��������g��"���O���)�)�_ @LM9�Dَ(�t���G���骼ʈ��&H"	A�wBI���P@I�4��,@l���v�77�1�h�J�u���42izs���Mx���Pױ3?qw$S�	�m�p